Title "CW Source check "

Osp Jobcontrol Verbosity=DEBUG  AllMon=0 AllMon=0

.option ingold=2 DELMAX=.1e-10 ACCURATE=1 RUNLVL=6 NUMDGT=8
.OPTION DCCAP=1 TNOM=27

.param PI=3.14159265358979
.param FourPI='4*3.1415926'
.param PIover2='3.1415926/2.0'
.param Noffset = 3.0e-4
%.param Non = '3.0  + Noffset'
%.param Noff = '3.012 + Noffset'

.param Noff = '1.6532'
.param Non = '1.6532'
.param NonWG = '1.4'

.param NMODES=1

* Voltage sources
v11 Mag1 0 DC = 1 
v12 Phi1 0 DC = 0

v21 Mag2 0 DC = 1 
v22 Phi2 0 DC = 0 

v31 Mag3 0 DC = 1 
v32 Phi3 0 DC = 0

v41 Mag4 0 DC = 1 
v42 Phi4 0 DC = 0 

v51 Mag5 0 DC = 1 
v52 Phi5 0 DC = 0

v3p51 Mag3p5 0 DC = 1 
v3p52 Phi3p5 0 DC = 0 

* lambda sweep Voltage
vcar vc 0 DC=1513

%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%

% circuit 5, One ring and 2 cross with waveguides

Osp CWSOURCE      Name = Rcw1 Nodes = [Mag1 Phi1 N11] MoName = CWmodel lambda = lam CarrierFreqNode=vc

Osp OpticalRing   Name = ring1 Nodes = [N11 N12 N13 N14] MoName = RingModel1


Osp WaveGuide  Name=wg1 Nodes = [N13 x11] MoName=WGmodel  
Osp WaveGuide  Name=wg2 Nodes = [N14 x12] MoName=WGmodel
  
Osp XCOUPLER    Name=wx1 Nodes = [x11 x12 x13 x14] MoName=WXmodel  

Osp WaveGuide  Name=wg3 Nodes = [x13 w3x1e] MoName=WGmodel  
Osp WaveGuide  Name=wg4 Nodes = [x14 w4x1n] MoName=WGmodel 


Osp XCOUPLER    Name=wx2 Nodes = [w3x1e x22 x23 x24] MoName=WXmodel

Osp WaveGuide  Name=wg5 Nodes = [x22 w2x2s] MoName=WGmodel
Osp WaveGuide  Name=wg6 Nodes = [x23 w3x2e] MoName=WGmodel  
Osp WaveGuide  Name=wg7 Nodes = [x24 w4x2n] MoName=WGmodel 

Osp MIRROR        Name = mirN12 Nodes = [N12] MoName = Mmodel
Osp MIRROR        Name = WGmir4x1n Nodes = [w4x1n] MoName = Mmodel 
Osp MIRROR        Name = WGmir2x2s Nodes = [w2x2s] MoName = Mmodel
Osp MIRROR        Name = WGmir3x2e Nodes = [w3x2e] MoName = Mmodel 
Osp MIRROR        Name = WGmir4x2n Nodes = [w4x2n] MoName = Mmodel
%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%

% Mirror Model
Osp Model Name = Mmodel   type = MIRROR Ref = 0.0 

% Source Model
Osp Model Name = CWmodel  type = CWSOURCE NumModes = NMODES lambda=lam



% Ring related Models  START

%Ring general Model statment
Osp Model Name = RingModel1 type = OptRing XC_model = XCmodel1 RingModel=RingFilter1 Radius = r1
Osp Model Name = RingModel2 type = OptRing XC_model = XCmodel1 RingModel=RingFilter1 Radius = r2
Osp Model Name = RingModel3 type = OptRing XC_model = XCmodel1 RingModel=RingFilter1 Radius = r3

% Coupling Model
Osp Model Name = XCmodel1  type = XCOUPLER Conjugate=0 c = C

% Filter model
Osp Model Name = RingFilter1 type = MultiLayerFilter FilterType=Explicit
+         N0=Non NF=Non TotalAtten = gain Index = [Non]  
  
% Ring related Models  END

% Xcouple model
Osp Model Name = WXmodel  type = XCOUPLER ElemType=WGUIDECROSS  NumModes = NMODES 
% +                         Through=0.9 Right=0.01 Left=0.01 Ref=0.1 



% WGuide model
Osp Model Name = WGmodel  type = WaveGuide  Length=1   neff=[Non]  N0=Non NF=Non
%Osp Model Name = WGmodel  type = WaveGuide  Length=1   neff=[NonWG]  N0=Non NF=Non

** gain is for pwr so sqrt is taken 
%.param gain='1'
.param gain='0.85'

.param r1='10.35'
.param r2='10.30'
.param r3='10.25'
.param C = '0.25'

.param lam=1513
.op 
.DC vcar 1510 1600 0.1
%.tran .1e-9 10e-9 nsolver=BACKE 

%.Monitor V Mag1 
%.Monitor V ring1 port=1 dir=IN


%.Monitor OptFields l5 Format=MagPhi Port=1 dir=IN  Pol=TE


% Outputs for circut 3.5, (ring1, x1, x1-4) // 20 outputs c2-
.Monitor OptPower ring1 Port=1 dir=IN Pol=TE  P0db=1 % C2
.Monitor OptPower ring1 Port=2 dir=IN Pol=TE  P0db=1 % C3
.Monitor OptPower ring1 Port=3 dir=IN Pol=TE  P0db=1 % C4
.Monitor OptPower ring1 Port=4 dir=IN Pol=TE  P0db=1 % C5

.Monitor OptPower ring1 Port=1 dir=OUT Pol=TE  P0db=1 % C6
.Monitor OptPower ring1 Port=2 dir=OUT Pol=TE  P0db=1 % C7
.Monitor OptPower ring1 Port=3 dir=OUT Pol=TE  P0db=1 % C8
.Monitor OptPower ring1 Port=4 dir=OUT Pol=TE  P0db=1 % C9

.Monitor OptPower wx1 Port=1 dir=IN Pol=TE  P0db=1 % C10
.Monitor OptPower wx1 Port=2 dir=IN Pol=TE  P0db=1 % C11
.Monitor OptPower wx1 Port=3 dir=IN Pol=TE  P0db=1 % C12
.Monitor OptPower wx1 Port=4 dir=IN Pol=TE  P0db=1 % C13

.Monitor OptPower wx1 Port=1 dir=OUT Pol=TE  P0db=1 % C14
.Monitor OptPower wx1 Port=2 dir=OUT Pol=TE  P0db=1 % C15
.Monitor OptPower wx1 Port=3 dir=OUT Pol=TE  P0db=1 % C16
.Monitor OptPower wx1 Port=4 dir=OUT Pol=TE  P0db=1 % C17

.Monitor OptPower wg4 Port=2 dir=IN Pol=TE  P0db=1 % C18
.Monitor OptPower wg4 Port=2 dir=OUT Pol=TE  P0db=1 % C19

.Monitor OptPower wx2 Port=1 dir=IN Pol=TE  P0db=1 % C20
.Monitor OptPower wx2 Port=2 dir=IN Pol=TE  P0db=1 % C21
.Monitor OptPower wx2 Port=3 dir=IN Pol=TE  P0db=1 % C22
.Monitor OptPower wx2 Port=4 dir=IN Pol=TE  P0db=1 % C23

.Monitor OptPower wx2 Port=1 dir=OUT Pol=TE  P0db=1 % C24
.Monitor OptPower wx2 Port=2 dir=OUT Pol=TE  P0db=1 % C25
.Monitor OptPower wx2 Port=3 dir=OUT Pol=TE  P0db=1 % C26
.Monitor OptPower wx2 Port=4 dir=OUT Pol=TE  P0db=1 % C27

.Monitor OptPower wg5 Port=2 dir=IN Pol=TE  P0db=1 % C28
.Monitor OptPower wg6 Port=2 dir=IN Pol=TE  P0db=1 % C29
.Monitor OptPower wg7 Port=2 dir=IN Pol=TE  P0db=1 % C30

.Monitor OptPower wg5 Port=2 dir=OUT Pol=TE  P0db=1 % C31
.Monitor OptPower wg6 Port=2 dir=OUT Pol=TE  P0db=1 % C32
.Monitor OptPower wg7 Port=2 dir=OUT Pol=TE  P0db=1 % C33

%.Monitor OptFields ring1 Format=MagPhi Port=1 dir=IN  Pol=TE %C22,23
%.Monitor OptFields ring1 Format=MagPhi Port=2 dir=IN  Pol=TE %C24,25
%.Monitor OptFields ring1 Format=MagPhi Port=3 dir=IN  Pol=TE %C26,27
%.Monitor OptFields ring1 Format=MagPhi Port=4 dir=IN  Pol=TE %C28,29

%.Monitor OptFields ring1 Format=MagPhi Port=1 dir=OUT  Pol=TE %C30,31
%.Monitor OptFields ring1 Format=MagPhi Port=2 dir=OUT  Pol=TE %C32,33
%.Monitor OptFields ring1 Format=MagPhi Port=3 dir=OUT  Pol=TE %C34,35
%.Monitor OptFields ring1 Format=MagPhi Port=4 dir=OUT  Pol=TE %C36,37

%.Monitor OptFields wx1 Format=MagPhi Port=1 dir=IN  Pol=TE %C38,39
%.Monitor OptFields wx1 Format=MagPhi Port=2 dir=IN  Pol=TE %C40,41
%.Monitor OptFields wx1 Format=MagPhi Port=3 dir=IN  Pol=TE %C42,43
%.Monitor OptFields wx1 Format=MagPhi Port=4 dir=IN  Pol=TE %C44,45

%.Monitor OptFields wx1 Format=MagPhi Port=1 dir=OUT  Pol=TE %C46,47
%.Monitor OptFields wx1 Format=MagPhi Port=2 dir=OUT  Pol=TE %C48,49
%.Monitor OptFields wx1 Format=MagPhi Port=3 dir=OUT  Pol=TE %C50,51
%.Monitor OptFields wx1 Format=MagPhi Port=4 dir=OUT  Pol=TE %C52,53


%.Monitor OptFields wg4 Format=MagPhi Port=2 dir=IN  Pol=TE %C56,57
%.Monitor OptFields wg4 Format=MagPhi Port=2 dir=Out  Pol=TE %C60,61

.end
